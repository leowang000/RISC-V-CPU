`include "global_params.v"

module reservation_station (
    input wire clk,
    input wire flush,
    
);
    
endmodule