`include "global_params.v"

module icache (
    
);
    
endmodule